module testbench;

endmodule : testbench